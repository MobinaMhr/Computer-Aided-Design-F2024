library verilog;
use verilog.vl_types.all;
entity Maxnet_NN_tb is
end Maxnet_NN_tb;
