library verilog;
use verilog.vl_types.all;
entity \Buffer\ is
    port(
        W0              : out    vl_logic_vector(31 downto 0);
        W1              : out    vl_logic_vector(31 downto 0);
        W2              : out    vl_logic_vector(31 downto 0);
        W3              : out    vl_logic_vector(31 downto 0);
        W4              : out    vl_logic_vector(31 downto 0);
        W5              : out    vl_logic_vector(31 downto 0);
        W6              : out    vl_logic_vector(31 downto 0);
        W7              : out    vl_logic_vector(31 downto 0);
        W8              : out    vl_logic_vector(31 downto 0);
        W9              : out    vl_logic_vector(31 downto 0);
        W10             : out    vl_logic_vector(31 downto 0);
        W11             : out    vl_logic_vector(31 downto 0);
        W12             : out    vl_logic_vector(31 downto 0);
        W13             : out    vl_logic_vector(31 downto 0);
        W14             : out    vl_logic_vector(31 downto 0);
        W15             : out    vl_logic_vector(31 downto 0)
    );
end \Buffer\;
